module alu_controller();
    
endmodule
